`timescale 1 ns / 1 ps
module SPI_0	
	#(
	parameter [5:0]  SPCRn_Address    = 6'h2C,  // I/O address for SPCR
	parameter [5:0]  SPSRn_Address    = 6'h2D,  // I/O address for SPSR
	parameter [5:0]  SPDRn_Address    = 6'h2E,  // I/O address for SPDR
	parameter [5:0]  SpiIRQ_Address   = 6'h11,
	// Memory interface addresses
	parameter [11:0] SPCRn_mem_Address  = 12'h04C,
	parameter [11:0] SPSRn_mem_Address  = 12'h04D,
	parameter [11:0] SPDRn_mem_Address  = 12'h04E
	)
	( 
	input             ireset,
	input             cp2,
	input [5:0]       IO_Addr,      // I/O bus address
	input             iore,
	input             iowe,
	output reg        out_en,
	input [7:0]       dbus_in,
	output reg [7:0]  dbus_out,
	// NVM part
	input             NVM_iore,
	input             NVM_iowe,
	input             SpiCRn,
	input             SpiSRn,
	input             SpiDRn,
	input logic       Disable_ireset,
	output logic [7:0] NVM_dbus_out,
	//
	input wire        miso_i,     // Master mode
	input wire        mosi_i,     // Slave mode
	input wire        sck_i,      // Slave mode
	input wire        ss_i,       // Slave/Master mode
	output wire       ss_o,       // Master mode
	output reg        miso_o,     // Slave mode
	output reg        mosi_o,     // Master mode
	output reg        sck_o,      // Master mode
	// IRQ
	output wire       SpiIRQ,
	input [5:0]       irqack_addr,
	input             irqack,
	// MEMORY INTERFACE PORTS added for RAM access:
	input [11:0]      ram_Addr,
	input             ramwe,
	input             ramre,
	// remaining I/O ports
	output          SPE0,
	output          MSTR0
	);
	reg [1:0] SpiAdr; //Adding
	assign SpiAdr = (SpiCRn) ? 2'b01 : 
					(SpiDRn) ? 2'b10 : 
					(SpiSRn) ? 2'b11 : 2'b00;
	reg [7:0]	SPCRn ;
	reg [7:0]	SPSRn ;
	// reg [7:0]	SPDRn ;
	// reg [7:0]	SPDRn_buf ;	

	reg SPIF_Next;
	reg WCOL_Next; 

	reg [7:0]           SPDR_Rc;
	reg [7:0]           SPDR_Rc_Next;
	reg [7:0]           SPDR_Sh_Current;
	reg [7:0]           SPDR_Sh_Next;
   
	reg [5:0]           Div_Next;
	reg [5:0]           Div_Current;
	reg                 Div_Toggle;
   
	reg                 DivCntMsb_Current;
	reg                 DivCntMsb_Next;
   
	localparam [3:0]     MstSMSt_Type_MstSt_Idle = 0,
						MstSMSt_Type_MstSt_B0 = 1,
						MstSMSt_Type_MstSt_B1 = 2,
						MstSMSt_Type_MstSt_B2 = 3,
						MstSMSt_Type_MstSt_B3 = 4,
						MstSMSt_Type_MstSt_B4 = 5,
						MstSMSt_Type_MstSt_B5 = 6,
						MstSMSt_Type_MstSt_B6 = 7,
						MstSMSt_Type_MstSt_B7 = 8;
	reg [3:0]           MstSMSt_Current;
	reg [3:0]           MstSMSt_Current_2;
	reg [3:0]           MstSMSt_Next;
   
	wire                TrStart;
   
	reg                 scko_Next;
	reg                 scko_Current;		//!!!
   
	reg                 UpdRcDataRg_Current;
	reg                 UpdRcDataRg_Next;
   
	reg                 TmpIn_Current;
	reg                 TmpIn_Next;
   
	// Slave
	reg                 sck_EdgeDetDFF;
	wire                SlvSampleSt;
   
	wire                SlvSMChangeSt;
   
	localparam [3:0]     SlvSMSt_Type_SlvSt_Idle = 0,
						SlvSMSt_Type_SlvSt_B0I = 1,
						SlvSMSt_Type_SlvSt_B0 = 2,
						SlvSMSt_Type_SlvSt_B1 = 3,
						SlvSMSt_Type_SlvSt_B2 = 4,
						SlvSMSt_Type_SlvSt_B3 = 5,
						SlvSMSt_Type_SlvSt_B4 = 6,
						SlvSMSt_Type_SlvSt_B5 = 7,
						SlvSMSt_Type_SlvSt_B6 = 8,
						SlvSMSt_Type_SlvSt_B6W = 9;
	reg [3:0]           SlvSMSt_Current;
	reg [3:0]           SlvSMSt_Next;
   
	// SIF clear SM
	reg                 SPIFClrSt_Current;
	reg                 SPIFClrSt_Next;
   
	// WCOL clear SM
	reg                 WCOLClrSt_Current;
	reg                 WCOLClrSt_Next;
   
	reg                 MstDSamp_Next;
	reg                 MstDSamp_Current;

	wire				SpiIRQ_Ack;
	reg					irst; //Adding
	assign	irst = ireset | Disable_ireset; //Adding
	function[7:0] Fn_RevBitVector;
		input [7:0]        InVector;
		input  integer    Dummy_Agr;
		begin
			Fn_RevBitVector = {InVector[0],InVector[1],InVector[2],InVector[3],InVector[4],InVector[5],InVector[6],InVector[7]};
		end
	endfunction

	assign SPE0 = SPCRn[6];
	assign MSTR0 = SPCRn[4];
	assign SpiIRQ_Ack = (irqack_addr == SpiIRQ_Address) && irqack ;
	
	always @(negedge irst or posedge cp2)
    begin : SPCRn_REG
        if (!irst) begin		// Reset
            SPCRn <= {8{1'b0}};
        end else begin		// Clock
            // Update on I/O access or RAM access
            if (((IO_Addr == SPCRn_Address) && iowe) ||
                ((ram_Addr == SPCRn_mem_Address) && ramwe)) begin
                SPCRn[7:5] <= dbus_in[7:5];
                SPCRn[3:0] <= dbus_in[3:0];
            end
            else if ( SpiCRn == 1 && NVM_iowe ) begin
                SPCRn[7:5] <= dbus_in[7:5];
                SPCRn[3:0] <= dbus_in[3:0];
            end
            case (SPCRn[4])
                1'b0 :
                    if ((IO_Addr == SPCRn_Address && iowe == 1'b1 && dbus_in[4] == 1'b1) ||
                        (ram_Addr == SPCRn_mem_Address && ramwe == 1'b1 && dbus_in[4] == 1'b1)) begin		
                        SPCRn[4] <= 1'b1;
                    end else if (SpiCRn == 1 && NVM_iowe && dbus_in[4] == 1'b1) begin
                        SPCRn[4] <= 1'b1;
                    end
                1'b1 :
                    if (((IO_Addr == SPCRn_Address && iowe == 1'b1 && dbus_in[4] == 1'b0) ||
                         (ram_Addr == SPCRn_mem_Address && ramwe == 1'b1 && dbus_in[4] == 1'b0)) || (ss_i == 1'b0)) begin 
                        SPCRn[4] <= 1'b0;
                    end else if ((SpiCRn == 1 && NVM_iowe && dbus_in[4] == 1'b0) || (ss_i == 1'b0)) begin
                        SPCRn[4] <= 1'b0;
                    end
            endcase
        end
    end
	
	always @(negedge irst or posedge cp2)
    begin : SPI2X_bit
        if (!irst) begin		// Reset
            SPSRn[0] <= 1'b0 ;
        end else begin		// Clock
            if (((IO_Addr == SPSRn_Address) && iowe) || ((ram_Addr == SPSRn_mem_Address) && ramwe) ||
                ((SpiSRn == 1) && (NVM_iowe == 1))) begin
                SPSRn[0] <= dbus_in[0];
            end
        end
    end
	
	always @(negedge irst or posedge cp2)
	begin : SeqPrc
		if (!irst) begin		// Reset
			SPSRn[7:1] <= {7{1'b0}};
			
			Div_Current <= {6{1'b0}};
			DivCntMsb_Current <= 1'b0;

			MstSMSt_Current <= MstSMSt_Type_MstSt_Idle;
			MstSMSt_Current_2 <= MstSMSt_Type_MstSt_Idle;
			SlvSMSt_Current <= SlvSMSt_Type_SlvSt_Idle;

			SPDR_Sh_Current <= {8{1'b1}};
			SPDR_Rc <= {8{1'b0}};

			sck_EdgeDetDFF <= 1'b0;
			SPIFClrSt_Current <= 1'b0;
			WCOLClrSt_Current <= 1'b0;

			sck_o <= 1'b0;
			scko_Current <= 1'b0;
			miso_o <= 1'b0;
			mosi_o <= 1'b0;

			TmpIn_Current <= 1'b0;
			UpdRcDataRg_Current <= 1'b0;
			MstDSamp_Current <= 1'b0;
		end else begin // Clock
			SPSRn[7] <= SPIF_Next;
			SPSRn[6] <= WCOL_Next;

			Div_Current <= Div_Next;
			DivCntMsb_Current <= DivCntMsb_Next;

			MstSMSt_Current <= MstSMSt_Next;
			MstSMSt_Current_2 <= MstSMSt_Next;

			SlvSMSt_Current <= SlvSMSt_Next;
			SPDR_Sh_Current <= SPDR_Sh_Next;
			SPDR_Rc <= SPDR_Rc_Next;
			sck_EdgeDetDFF <= sck_i;
			SPIFClrSt_Current <= SPIFClrSt_Next;
			WCOLClrSt_Current <= WCOLClrSt_Next;

			scko_Current <= scko_Next;
			sck_o <= scko_Next;
			miso_o <= SPDR_Sh_Next[7];
			mosi_o <= SPDR_Sh_Next[7];

			TmpIn_Current <= TmpIn_Next;
			UpdRcDataRg_Current <= UpdRcDataRg_Next;
			MstDSamp_Current <= MstDSamp_Next;
		end
	end // SeqPrc 
	
	// always @(MstSMSt_Current or Div_Current or SPCRn or SPSRn)
	always_comb
	begin : DividerToggleComb
		Div_Toggle = 1'b0;
		if (MstSMSt_Current != MstSMSt_Type_MstSt_Idle) begin
			if (SPSRn[0] == 1'b1) begin		// Extended mode
				case (SPCRn[1:0])
					2'b00 :		// fosc /2
						if (Div_Current == 6'b000000) begin
							Div_Toggle = 1'b1;
						end
					2'b01 :		// fosc /8
						if (Div_Current == 6'b000011) begin
							Div_Toggle = 1'b1;
						end
					2'b10 :		// fosc /32
						if (Div_Current == 6'b001111) begin
							Div_Toggle = 1'b1;
						end
					2'b11 :		// fosc /64
						if (Div_Current == 6'b011111) begin
							Div_Toggle = 1'b1;
						end
					// default :
					// 	Div_Toggle = 1'b0;
				endcase
			end else begin // Normal mode
				case (SPCRn[1:0])
					2'b00 :		// fosc /4	  
						if (Div_Current == 6'b000001) begin
							Div_Toggle = 1'b1;
						end
					2'b01 :		// fosc /16
						if (Div_Current == 6'b000111) begin
							Div_Toggle = 1'b1;
						end
					2'b10 :		// fosc /64
						if (Div_Current == 6'b011111) begin
							Div_Toggle = 1'b1;
						end
					2'b11 :		// fosc /128
						if (Div_Current == 6'b111111) begin
							Div_Toggle = 1'b1;
						end
					// default :
					// 	Div_Toggle = 1'b0;
				endcase
			end
		end
	end
   
	// always @(MstSMSt_Current_2 or Div_Current or DivCntMsb_Current or Div_Toggle)
	always_comb
	begin : DividerNextComb
		Div_Next = Div_Current;
		DivCntMsb_Next = DivCntMsb_Current;
		if (MstSMSt_Current != MstSMSt_Type_MstSt_Idle) begin
			if (Div_Toggle == 1'b1)begin
				Div_Next = {6{1'b0}};
				DivCntMsb_Next = (~DivCntMsb_Current);
			end else begin
				Div_Next = Div_Current + 1;
			end
		end
    end

	// always @(MstSMSt_Current or Div_Current or DivCntMsb_Current or Div_Toggle)
	// begin : DividerNextComb
	// 	case (MstSMSt_Current)
	// 		MstSMSt_Type_MstSt_Idle : begin
	// 			Div_Next = Div_Current;
	// 			DivCntMsb_Next = DivCntMsb_Current; 
	// 			end
	// 		default: 
	// 			if (Div_Toggle == 1'b1)begin
	// 				Div_Next = {6{1'b0}};
	// 				DivCntMsb_Next = (~DivCntMsb_Current);
	// 			end else begin
	// 				Div_Next = Div_Current + 1;
	// 				DivCntMsb_Next = DivCntMsb_Current;
	// 			end
	// 	endcase
    // end
   
	assign TrStart = ((IO_Addr == SPDRn_Address & iowe == 1'b1 & SPCRn[6] == 1'b1) | 
	                 (ram_Addr == SPDRn_mem_Address & ramwe == 1'b1 & SPCRn[6] == 1'b1) |
	                 (SpiDRn == 1 & NVM_iowe == 1'b1 & SPCRn[6] == 1'b1)) ? 1'b1 : 1'b0;
   
   // Transmitter Master Mode Shift Control SM
   
	// always @(MstSMSt_Current or DivCntMsb_Current or Div_Toggle or TrStart or SPCRn)
	always_comb
	begin : MstSmNextComb
		MstSMSt_Next = MstSMSt_Current;
		case (MstSMSt_Current)
			MstSMSt_Type_MstSt_Idle :
				if (TrStart == 1'b1 & SPCRn[4] == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B0;
				end
			MstSMSt_Type_MstSt_B0 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B1;
				end
			MstSMSt_Type_MstSt_B1 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B2;
				end
			MstSMSt_Type_MstSt_B2 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B3;
				end
			MstSMSt_Type_MstSt_B3 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B4;
				end
			MstSMSt_Type_MstSt_B4 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B5;
				end
			MstSMSt_Type_MstSt_B5 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B6;
				end
			MstSMSt_Type_MstSt_B6 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_B7;
				end
			MstSMSt_Type_MstSt_B7 :
				if (DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) begin
					MstSMSt_Next = MstSMSt_Type_MstSt_Idle;
				end
			// default :
			// 	MstSMSt_Next = MstSMSt_Type_MstSt_Idle;
		endcase
	end
   
   
	always_comb
	begin : SPIFClrCombProc
		SPIFClrSt_Next = SPIFClrSt_Current;
		case (SPIFClrSt_Current)
			1'b0 :
				if ((((IO_Addr == SPSRn_Address & iore == 1'b1) | 
				     (ram_Addr == SPSRn_mem_Address & ramre == 1'b1) |
				     (SpiSRn == 1 & NVM_iore == 1'b1)) & 
				     SPSRn[7] == 1'b1 & SPCRn[6] == 1'b1)) begin
					SPIFClrSt_Next = 1'b1;
				end
			1'b1 :
				if (((IO_Addr == SPDRn_Address & (iore == 1'b1 | iowe == 1'b1)) | 
				    (ram_Addr == SPDRn_mem_Address & (ramre == 1'b1 | ramwe == 1'b1)) |
				    (SpiDRn == 1 & (NVM_iowe == 1 | NVM_iore == 1'b1)))) begin
					SPIFClrSt_Next = 1'b0;
				end
		endcase
	end  //SPIFClrCombProc
      
      
    always_comb
    begin : WCOLClrCombProc
        WCOLClrSt_Next = WCOLClrSt_Current;
        case (WCOLClrSt_Current)
			1'b0 :
				if ((((IO_Addr == SPSRn_Address & iore == 1'b1) |
				     (ram_Addr == SPSRn_mem_Address & ramre == 1'b1) |
				     (SpiSRn == 1 & NVM_iore == 1'b1)) & 
				     SPSRn[6] == 1'b1)) begin 
					WCOLClrSt_Next = 1'b1;
				end
            1'b1 :
				if (((IO_Addr == SPDRn_Address & (iore == 1'b1 | iowe == 1'b1)) |
				    (ram_Addr == SPDRn_mem_Address & (ramre == 1'b1 | ramwe == 1'b1)) |
				    (SpiDRn == 1 & (NVM_iowe == 1'b1 | NVM_iore == 1'b1)))) begin
					WCOLClrSt_Next = 1'b0;
				end
            default :
				WCOLClrSt_Next = WCOLClrSt_Current;
        endcase
    end //WCOLClrCombProc
         
         
    always_comb
    begin : MstDataSamplingComb
        MstDSamp_Next = 1'b0;
        case (MstDSamp_Current)
            1'b0 :
				if (MstSMSt_Current != MstSMSt_Type_MstSt_Idle) begin
                    if (SPCRn[2] == SPCRn[3]) begin
                        if (scko_Next == 1'b1 & scko_Current == 1'b0) begin		// Rising edge 	  
                           MstDSamp_Next = 1'b1;
						end
                    end else begin // CPHA/=CPOL
                        if (scko_Next == 1'b0 & scko_Current == 1'b1) begin		// Falling edge 	  
                           MstDSamp_Next = 1'b1;
						end
					end
                end
            1'b1 :
                MstDSamp_Next = 1'b0;
            // default :
            //     MstDSamp_Next = 1'b0;
        endcase
    end // MstDataSamplingComb
            
            //
            
    always_comb
    begin : DRLatchComb
        UpdRcDataRg_Next = 1'b0;
        case (UpdRcDataRg_Current)
            1'b0 :
                if ((SPCRn[4] == 1'b1 & MstSMSt_Current != MstSMSt_Type_MstSt_Idle & MstSMSt_Next == MstSMSt_Type_MstSt_Idle) | (SPCRn[4] == 1'b0 & SlvSMSt_Current != SlvSMSt_Type_SlvSt_Idle & SlvSMSt_Next == SlvSMSt_Type_SlvSt_Idle)) begin
                    UpdRcDataRg_Next = 1'b1;
				end
            1'b1 :
                UpdRcDataRg_Next = 1'b0;
			// default :
			// 	UpdRcDataRg_Next = 1'b0;
        endcase
    end
            
            
    always_comb
    begin : TmpInComb
        TmpIn_Next = TmpIn_Current;
        if (SPCRn[4] == 1'b1 & MstDSamp_Current == 1'b1) begin		// Master mode
            TmpIn_Next = miso_i;
        end else if (SPCRn[4] == 1'b0 & SlvSampleSt == 1'b1 & ss_i == 1'b0) begin		// Slave mode ???
            TmpIn_Next = mosi_i;
		end
    end

    always_comb
    begin : ShiftRgComb
        SPDR_Sh_Next = SPDR_Sh_Current;
        if (TrStart == 1'b1 & (MstSMSt_Current == MstSMSt_Type_MstSt_Idle & SlvSMSt_Current == SlvSMSt_Type_SlvSt_Idle & (~(SPCRn[4] == 1'b0 & SlvSampleSt == 1'b1 & ss_i == 1'b0)))) begin		// Load
            if (SPCRn[5] == 1'b1) begin		// the LSB of the data word is transmitted first
				SPDR_Sh_Next = Fn_RevBitVector(dbus_in, 8);
            end else begin// the MSB of the data word is transmitted first
                SPDR_Sh_Next = dbus_in;
			end
        end else if (SPCRn[4] == 1'b1 & UpdRcDataRg_Current == 1'b1) begin	 	// ???
                  SPDR_Sh_Next[7] = 1'b1;
        end else if ((SPCRn[4] == 1'b1 & MstSMSt_Current != MstSMSt_Type_MstSt_Idle & DivCntMsb_Current == 1'b1 & Div_Toggle == 1'b1) | (SPCRn[4] == 1'b0 & SlvSMSt_Current != SlvSMSt_Type_SlvSt_Idle & SlvSMChangeSt == 1'b1 & ss_i == 1'b0)) begin
                  // Shift
            SPDR_Sh_Next = {SPDR_Sh_Current[7 - 1:0], TmpIn_Current};
		end
	end //ShiftRgComb
               
               
	always_comb
	begin : sckoGenComb
		scko_Next = scko_Current;
		if ((IO_Addr == SPCRn_Address & iowe == 1'b1) || 
		    (ram_Addr == SPCRn_mem_Address & ramwe == 1'b1)) begin  // Write to SPCR
			scko_Next = dbus_in[3];		// CPOL
		end else if (TrStart == 1'b1 & SPCRn[2] == 1'b1 & MstSMSt_Current == MstSMSt_Type_MstSt_Idle) begin
			scko_Next = (~SPCRn[3]);
		end else if (MstSMSt_Current != MstSMSt_Type_MstSt_Idle & MstSMSt_Next == MstSMSt_Type_MstSt_Idle) begin		// "Parking"
			scko_Next = SPCRn[3];
		end else if (MstSMSt_Current != MstSMSt_Type_MstSt_Idle & DivCntMsb_Current != DivCntMsb_Next) begin
			scko_Next = (~scko_Current);
		end
	end
               
    // Receiver data register
               
	always_comb
	begin : SPDRRcComb
		SPDR_Rc_Next = SPDR_Rc;
		if (UpdRcDataRg_Current == 1'b1) begin
			if (SPCRn[4] == 1'b0 & SPCRn[2] == 1'b1) begin
				if (SPCRn[5] == 1'b1) begin		// the LSB of the data word is transmitted first
					SPDR_Rc_Next = Fn_RevBitVector({SPDR_Sh_Current[7 - 1:0], TmpIn_Current}, 2);
				end else begin // the MSB of the data word is transmitted first
					SPDR_Rc_Next = {SPDR_Sh_Current[7 - 1:0], TmpIn_Current};
				end
			end else begin
				if (SPCRn[5] == 1'b1) begin		// the LSB of the data word is transmitted first
					SPDR_Rc_Next = Fn_RevBitVector(SPDR_Sh_Current, 8);
				end else begin // the MSB of the data word is transmitted first
					SPDR_Rc_Next = SPDR_Sh_Current;
				end
			end
		end
	end
               
	//****************************************************************************************			
	// Slave
	//****************************************************************************************

	// Rising edge 
	assign SlvSampleSt = (((sck_EdgeDetDFF == 1'b0 & sck_i == 1'b1 & SPCRn[3] == SPCRn[2]) | (sck_EdgeDetDFF == 1'b1 & sck_i == 1'b0 & SPCRn[3] != SPCRn[2]))) ? 1'b1 : 		// Falling edge
						1'b0;

	// Falling edge 
	assign SlvSMChangeSt = (((sck_EdgeDetDFF == 1'b1 & sck_i == 1'b0 & SPCRn[3] == SPCRn[2]) | (sck_EdgeDetDFF == 1'b0 & sck_i == 1'b1 & SPCRn[3] != SPCRn[2]))) ? 1'b1 : 		// Rising edge
						  1'b0;

	// Slave Master Mode Shift Control SM
               
	always_comb
	begin : SlvSMNextComb
		SlvSMSt_Next = SlvSMSt_Current;
		if (ss_i == 1'b0) begin
			case (SlvSMSt_Current)
				SlvSMSt_Type_SlvSt_Idle :
					if (SPCRn[4] == 1'b0) begin
						if (SPCRn[2] == 1'b1) begin
							if (SlvSMChangeSt == 1'b1) begin
								SlvSMSt_Next = SlvSMSt_Type_SlvSt_B0;
							end
						end else begin //	CPHA='0'
							if (SlvSampleSt == 1'b1) begin
								SlvSMSt_Next = SlvSMSt_Type_SlvSt_B0I;
							end
						end
					end
				SlvSMSt_Type_SlvSt_B0I :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B0;
					end
				SlvSMSt_Type_SlvSt_B0 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B1;
					end
				SlvSMSt_Type_SlvSt_B1 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B2;
					end
				SlvSMSt_Type_SlvSt_B2 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B3;
					end
				SlvSMSt_Type_SlvSt_B3 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B4;
					end
				SlvSMSt_Type_SlvSt_B4 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B5;
					end
				SlvSMSt_Type_SlvSt_B5 :
					if (SlvSMChangeSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_B6;
					end
				SlvSMSt_Type_SlvSt_B6 :
					if (SlvSMChangeSt == 1'b1) begin
						if (SPCRn[2] == 1'b0) begin
							SlvSMSt_Next = SlvSMSt_Type_SlvSt_Idle;
						end else begin// CPHA='1'
							SlvSMSt_Next = SlvSMSt_Type_SlvSt_B6W;
						end
					end
				SlvSMSt_Type_SlvSt_B6W :
					if (SlvSampleSt == 1'b1) begin
						SlvSMSt_Next = SlvSMSt_Type_SlvSt_Idle;
					end
				default :
					SlvSMSt_Next = SlvSMSt_Type_SlvSt_Idle;
			endcase
		end
	end
               
               
	// always @(adr or iowe or dbus_in or ss_b_resync or SPCR)
	// begin: MSTRGenComb
		// MSTR_Next = `MSTR;
		// case (`MSTR)
			// 1'b0 :
				// if (adr == SPCR_Address & iowe == 1'b1 & dbus_in[4] == 1'b1)		// TBD (ss_b_resync='0')
					// MSTR_Next = 1'b1;
			// 1'b1 :
				// if ((adr == SPCR_Address & iowe == 1'b1 & dbus_in[4] == 1'b0) | (ss_b_resync == 1'b0))
					// MSTR_Next = 1'b0;
			// default :
				// MSTR_Next = `MSTR;
		// endcase
	// end


	always_comb
	begin : WCOLGenComb
		WCOL_Next = SPSRn[6];
		case (SPSRn[6])
			1'b0 :
				if ((((IO_Addr == SPDRn_Address & iowe == 1'b1) | 
				     (ram_Addr == SPDRn_mem_Address & ramwe == 1'b1) |
				     (SpiDRn == 1 & NVM_iowe == 1)) & 
				     ((SPCRn[4] == 1'b0 & (SlvSMSt_Current != SlvSMSt_Type_SlvSt_Idle | (SlvSampleSt == 1'b1 & ss_i == 1'b0))) | 
				     (SPCRn[4] == 1'b1 & MstSMSt_Current != MstSMSt_Type_MstSt_Idle))))
					WCOL_Next = 1'b1;
			1'b1 :
				if (((((IO_Addr == SPDRn_Address & (iowe == 1'b1 | iore == 1'b1)) |
				      (ram_Addr == SPDRn_mem_Address & (ramwe == 1'b1 | ramre == 1'b1)) |
				      (SpiDRn == 1 & (NVM_iowe == 1 | NVM_iore == 1))) & WCOLClrSt_Current == 1'b1) & 
				      (~(((IO_Addr == SPDRn_Address & iowe == 1'b1) |
				         (ram_Addr == SPDRn_mem_Address & ramwe == 1'b1) |
				         (SpiDRn == 1 & NVM_iowe == 1)) & 
				         ((SPCRn[4] == 1'b0 & (SlvSMSt_Current != SlvSMSt_Type_SlvSt_Idle | (SlvSampleSt == 1'b1 & ss_i == 1'b0))) | 
				         (SPCRn[4] == 1'b1 & MstSMSt_Current != MstSMSt_Type_MstSt_Idle))))))
					WCOL_Next = 1'b0;
		endcase
	end


	always_comb
	begin : SPIFGenComb
		SPIF_Next = SPSRn[7];
		case (SPSRn[7])
			1'b0 :
				if ((SPCRn[4] == 1'b0 & SlvSMSt_Current != SlvSMSt_Type_SlvSt_Idle & SlvSMSt_Next == SlvSMSt_Type_SlvSt_Idle) | 
				   (SPCRn[4] == 1'b1 & MstSMSt_Current != MstSMSt_Type_MstSt_Idle & MstSMSt_Next == MstSMSt_Type_MstSt_Idle)| (SPCRn[4] == 1'b1 & ss_i == 1'b0))
					SPIF_Next = 1'b1;
			1'b1 :
				if (((((IO_Addr == SPDRn_Address & (iowe == 1'b1 | iore == 1'b1)) | 
				      (ram_Addr == SPDRn_mem_Address & (ramwe == 1'b1 | ramre == 1'b1)) |
				      (SpiDRn == 1 & (NVM_iore == 1 | NVM_iowe == 1))) & SPIFClrSt_Current == 1'b1) | 
				      SpiIRQ_Ack == 1'b1))
					SPIF_Next = 1'b0;
		endcase
	end

	//*************************************************************************************

	// IRQ
	assign SpiIRQ = SPCRn[7] & SPSRn[7];
	
	always @(*)
    begin: OutMuxComb

        if (ramre) begin
            case (ram_Addr)
                SPCRn_mem_Address: begin
                    dbus_out <= SPCRn;
                    out_en <= 1'b1;
                end
                SPSRn_mem_Address: begin
                    dbus_out <= SPSRn;
                    out_en <= 1'b1;
                end
                SPDRn_mem_Address: begin
                    dbus_out <= SPDR_Rc;
                    out_en <= 1'b1;
                end
                default: begin
                    dbus_out <= {8{1'b0}};
                    out_en <= 1'b0;
                end
            endcase
        end else begin
            case (IO_Addr)
                SPCRn_Address: begin
                    dbus_out <= SPCRn;
                    out_en <= iore;
                end
                SPSRn_Address: begin
                    dbus_out <= SPSRn;
                    out_en <= iore;
                end
                SPDRn_Address: begin
                    dbus_out <= SPDR_Rc;
                    out_en <= iore;
                end
                default: begin
                    dbus_out <= {8{1'b0}};
                    out_en <= 1'b0;
                end
            endcase
        end
    end

endmodule